netcdf OCEAN_SURFACE_FRESHWATER_FLUXES_mon_mean_1992-02_ECCO_V4r4_latlon_0p50deg {
dimensions:
	time = 1 ;
	latitude = 360 ;
	longitude = 720 ;
	nv = 2 ;
variables:
	int time(time) ;
		time:axis = "T" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "center time of averaging period or time of snapshot" ;
		time:standard_name = "time" ;
		time:units = "days since 1992-02-15 12:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:comment = "uniform grid spacing from -89.75 to 89.75 by 0.5" ;
		latitude:coverage_content_type = "coordinate" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:comment = "uniform grid spacing from -179.75 to 179.75 by 0.5" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	int time_step(time) ;
		time_step:coverage_content_type = "coordinate" ;
		time_step:long_name = "model time step [hours since 1992-01-01T12:00:00" ;
		time_step:units = "hours" ;
	float EXFpreci(time, latitude, longitude) ;
		EXFpreci:_FillValue = 9.96921e+36f ;
		EXFpreci:comment = "Precipitation rate. Note: sum of ERA-Interim precipitation and the control adjustment." ;
		EXFpreci:coverage_content_type = "modelResult" ;
		EXFpreci:direction = ">0 increases salinity (SALT)" ;
		EXFpreci:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE; FRESH WATER FLUX; PRECIPITATION; PRECIPITATION RATE; TOTAL SURFACE PRECIPITATION RATE" ;
		EXFpreci:long_name = "Precipitation rate" ;
		EXFpreci:standard_name = "lwe_precipitation_rate" ;
		EXFpreci:units = "m s-1" ;
		EXFpreci:coordinates = "time latitude longitude time_step" ;
	float latitude_bnds(latitude, nv) ;
		latitude_bnds:coverage_content_type = "coordinate" ;
		latitude_bnds:long_name = "latitude bounds of lat-lon grid cells" ;
	float longitude_bnds(longitude, nv) ;
		longitude_bnds:coverage_content_type = "coordinate" ;
		longitude_bnds:long_name = "longitude bounds of lat-lon grid cells" ;
	int time_bnds(time, nv) ;
		time_bnds:coverage_content_type = "coordinate" ;
		time_bnds:long_name = "start and stop time of period or time of snapshot" ;
		time_bnds:units = "days since 1992-02-01 00:00:00" ;
		time_bnds:calendar = "proleptic_gregorian" ;
	float EXFevap(time, latitude, longitude) ;
		EXFevap:_FillValue = 9.96921e+36f ;
		EXFevap:comment = "Open ocean evaporation. Note: calculated using the bulk formula following Large and Yeager, 2004, NCAR/TN-460+STR." ;
		EXFevap:coverage_content_type = "modelResult" ;
		EXFevap:direction = ">0 increases salinity (SALT)" ;
		EXFevap:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE; EVAPORATION; FRESH WATER FLUX" ;
		EXFevap:long_name = "Evaporation rate" ;
		EXFevap:standard_name = "lwe_water_evaporation_rate" ;
		EXFevap:units = "m s-1" ;
		EXFevap:coordinates = "time latitude longitude time_step" ;
	float EXFroff(time, latitude, longitude) ;
		EXFroff:_FillValue = 9.96921e+36f ;
		EXFroff:comment = "River runoff freshwater flux. Note: not adjusted by the optimization." ;
		EXFroff:coverage_content_type = "modelResult" ;
		EXFroff:direction = ">0 increases salinity (SALT)" ;
		EXFroff:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE" ;
		EXFroff:long_name = "River runoff" ;
		EXFroff:standard_name = "surface_runoff_flux" ;
		EXFroff:units = "m s-1" ;
		EXFroff:coordinates = "time latitude longitude time_step" ;
	float SIsnPrcp(time, latitude, longitude) ;
		SIsnPrcp:_FillValue = 9.96921e+36f ;
		SIsnPrcp:comment = "Snow precipitation rate over sea-ice, averaged over the entire model grid cell.   . " ;
		SIsnPrcp:coverage_content_type = "modelResult" ;
		SIsnPrcp:direction = ">0 increases snow thickness (HSNOW)" ;
		SIsnPrcp:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SEA ICE; SNOW/ICE; FRESH WATER FLUX; PRECIPITATION; PRECIPITATION RATE" ;
		SIsnPrcp:long_name = "Snow precipitation on sea-ice" ;
		SIsnPrcp:standard_name = "snowfall_flux" ;
		SIsnPrcp:units = "kg m-2 s-1" ;
		SIsnPrcp:coordinates = "time latitude longitude time_step" ;
	float EXFempmr(time, latitude, longitude) ;
		EXFempmr:_FillValue = 9.96921e+36f ;
		EXFempmr:comment = "Net freshwater flux out of the liquid ocean from precipitation, evaporation, and runoff and excluding freshwater fluxes involving sea-ice and snow. Note: calculated as EXFevap-EXFpreci-EXFroff." ;
		EXFempmr:coverage_content_type = "modelResult" ;
		EXFempmr:direction = ">0 increases salinity (SALT)" ;
		EXFempmr:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE; EVAPORATION; FRESH WATER FLUX" ;
		EXFempmr:long_name = "Net freshwater flux out of the ocean from precipitation, evaporation, and runoff" ;
		EXFempmr:units = "m s-1" ;
		EXFempmr:coordinates = "time latitude longitude time_step" ;
	float oceFWflx(time, latitude, longitude) ;
		oceFWflx:_FillValue = 9.96921e+36f ;
		oceFWflx:comment = "Net freshwater flux into the ocean including contributions from runoff, evaporation, precipitation, and mass exchange with sea-ice due to melting and freezing and snow melting. Note: \'oceFWflx\' does NOT include freshwater fluxes between the atmosphere and sea-ice and snow. The variable \'SIatmFW\' accounts for freshwater fluxes out of the combined ocean+sea-ice+snow reservoir." ;
		oceFWflx:coverage_content_type = "modelResult" ;
		oceFWflx:direction = ">0 decreases salinity (SALT)" ;
		oceFWflx:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; ATMOSPHERE; FRESH WATER FLUX" ;
		oceFWflx:long_name = "Net freshwater flux into the ocean" ;
		oceFWflx:standard_name = "water_flux_into_sea_water" ;
		oceFWflx:units = "kg m-2 s-1" ;
		oceFWflx:coordinates = "time latitude longitude time_step" ;
	float SIatmFW(time, latitude, longitude) ;
		SIatmFW:_FillValue = 9.96921e+36f ;
		SIatmFW:comment = "Net freshwater flux into the combined liquid ocean, sea-ice, and snow reservoirs from the atmosphere and runoff.. Note: freshwater fluxes BETWEEN the liquid ocean and sea-ice or snow reservoirs do not contribute to SIatmFW.  SIatmFW counts all fluxes to/from the atmosphere that change the TOTAL freshwater stored in the combined liquid ocean, sea-ice, and snow reservoirs." ;
		SIatmFW:coverage_content_type = "modelResult" ;
		SIatmFW:direction = ">0 increases salinity (SALT)" ;
		SIatmFW:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SEA ICE; SNOW/ICE; FRESH WATER FLUX" ;
		SIatmFW:long_name = "Net freshwater flux into the open ocean, sea-ice, and snow" ;
		SIatmFW:standard_name = "surface_upward_water_flux" ;
		SIatmFW:units = "kg m-2 s-1" ;
		SIatmFW:coordinates = "time latitude longitude time_step" ;
	float SFLUX(time, latitude, longitude) ;
		SFLUX:_FillValue = 9.96921e+36f ;
		SFLUX:comment = "The rate of change of total ocean salinity due to freshwater fluxes across the liquid surface and the addition or removal of mass. Note:  the global area integral of \'SFLUX\'  matches the time-derivative of total ocean salinity (psu s-1).  Unlike \'oceFWflx\', \'SFLUX\' includes the contribution to the total ocean salinity from changing ocean mass (e.g. from the addition or removal of freshwater in \'oceFWflx\'). " ;
		SFLUX:coverage_content_type = "modelResult" ;
		SFLUX:direction = ">0 increases salinity (SALT)" ;
		SFLUX:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SALT TRANSPORT" ;
		SFLUX:long_name = "Rate of change of total ocean salinity per m2 accounting for mass fluxes." ;
		SFLUX:units = "g m-2 s-1" ;
		SFLUX:coordinates = "time latitude longitude time_step" ;
	float SIacSubl(time, latitude, longitude) ;
		SIacSubl:_FillValue = 9.96921e+36f ;
		SIacSubl:comment = "Freshwater flux to the atmosphere due to sublimation-deposition of snow or ice. Positive values imply sublimation from ice/snow to vapor, negative values imply deposition from atmospheric moisture" ;
		SIacSubl:coverage_content_type = "modelResult" ;
		SIacSubl:direction = ">0 decreases snow or sea-ice thickness (HSNOW or HEFF)" ;
		SIacSubl:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SEA ICE; SNOW/ICE" ;
		SIacSubl:long_name = "Freshwater flux to the atmosphere due to sublimation-deposition of snow or ice" ;
		SIacSubl:standard_name = "water_sublimation_flux" ;
		SIacSubl:units = "kg m-2 s-1" ;
		SIacSubl:coordinates = "time latitude longitude time_step" ;
	float SIrsSubl(time, latitude, longitude) ;
		SIrsSubl:_FillValue = 9.96921e+36f ;
		SIrsSubl:comment = "Residual freshwater flux by sublimation to remove water from or add water to ocean. When implied sublimation freshwater flux \'SIacSubl\' is larger than availabe sea-ice/snow, \'SIrsSubl\' is positive and water is removed from ocean. Note: freshwater flux by sublimation that is to remove water from the ocean when it is positive." ;
		SIrsSubl:coverage_content_type = "modelResult" ;
		SIrsSubl:direction = ">0 decreases ocean volume" ;
		SIrsSubl:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SEA ICE; SNOW/ICE; FRESH WATER FLUX" ;
		SIrsSubl:long_name = "Residual sublimation freshwater flux" ;
		SIrsSubl:units = "kg m-2 s-1" ;
		SIrsSubl:coordinates = "time latitude longitude time_step" ;
	float SIfwThru(time, latitude, longitude) ;
		SIfwThru:_FillValue = 9.96921e+36f ;
		SIfwThru:comment = "Precipitation over sea-ice covered regions reaching ocean through sea-ice. Note: Precipitation over sea-ice covered regions that directly reaches ocean through the sea-ice. It is not due to melt of sea-ice/snow." ;
		SIfwThru:coverage_content_type = "modelResult" ;
		SIfwThru:direction = ">0 increases ocean volume" ;
		SIfwThru:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE; OCEANS; SEA ICE; SNOW/ICE; FRESH WATER FLUX; PRECIPITATION; PRECIPITATION RATE; TOTAL SURFACE PRECIPITATION RATE" ;
		SIfwThru:long_name = "Precipitation through sea-ice" ;
		SIfwThru:units = "kg m-2 s-1" ;
		SIfwThru:coordinates = "time latitude longitude time_step" ;

// global attributes:
		:acknowledgement = "This research was carried out by the Jet Propulsion Laboratory, managed by the California Institute of Technology under a contract with the National Aeronautics and Space Administration." ;
		:author = "Ian Fenty and Ou Wang" ;
		:cdm_data_type = "Grid" ;
		:comment = "These fields are provided on a regular lat-lon grid. They have been mapped to the regular lat-lon grid from the original ECCO lat-lon-cap 90 (llc90) native model grid." ;
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:coordinates = "time latitude longitude time_step latitude_bnds longitude_bnds time_bnds" ;
		:creator_email = "ecco-group@mit.edu" ;
		:creator_institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:creator_name = "ECCO Consortium" ;
		:creator_type = "group" ;
		:creator_url = "https://ecco.jpl.nasa.gov" ;
		:date_created = "TBD_DATASET" ;
		:date_issued = "2020-09-02T15:35:07.574548" ;
		:date_metadata_modified = "2020-09-02T15:35:07.574545" ;
		:date_modified = "2020-09-02T15:35:07.574537" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 90. ;
		:geospatial_lat_min = -90. ;
		:geospatial_lat_resolution = 0.5 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 180. ;
		:geospatial_lon_min = -180. ;
		:geospatial_lon_resolution = 0.5 ;
		:geospatial_lon_units = "degrees_east" ;
		:grid_mapping_name = "latitude_longitude" ;
		:history = "Inaugural release of an ECCO \"Central Estimate\" solution to PO.DAAC" ;
		:id = "TBD_DOI" ;
		:institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:keywords = "ECCO, State Estimate, Estimating the Circulation and Climate of the Ocean" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "Public Domain" ;
		:naming_authority = "gov.nasa.jpl" ;
		:nx = 720 ;
		:ny = 360 ;
		:platform = "ERS-1/2, TOPEX/Poseidon, GFO, ENVISAT, Jason-1, Jason-2, CryoSat-2, SARAL/AltiKa, Jason-3, AVHRR, Aquarius, SSM/I, SSMIS, GRACE, DTU17MDT, Argo, WOCE, GO-SHIP, MEOP, ITP" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:processing_level = "L4" ;
		:product_name = "TBD_FILENAME" ;
		:product_time_coverage_end = "2017-12-31T12:00:00" ;
		:product_time_coverage_start = "1992-01-01T12:00:00" ;
		:product_version = "Version 4, Release 4" ;
		:program = "NASA Physical Oceanography, Cryosphere, Modeling, Analysis, and Prediction (MAP)" ;
		:project = "Estimating the Circulation and Climate of the Ocean (ECCO)" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_institution = "PO.DAAC" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center (PO.DAAC)" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:references = "ECCO Consortium, Fukumori, I., Wang, O., Fenty, I., Forget, G., Heimbach, P., & Ponte, R. M. 2020. Synopsis of the ECCO Central Production Global Ocean and Sea-Ice State Estimate (Version 4 Release 4).doi:10.5281/zenodo.3765929" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:summary = "ocean and sea-ice surface freshwater fluxes" ;
		:time_coverage_duration = "P1M" ;
		:time_coverage_end = "1992-03-01T00:00:00.000000000" ;
		:time_coverage_resolution = "P1M" ;
		:time_coverage_start = "1992-02-01T00:00:00.000000000" ;
		:title = "ocean and sea-ice surface freshwater fluxes" ;
		:uuid = "TBD_DATASET" ;
}
