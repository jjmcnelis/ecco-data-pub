netcdf OCEAN_PRES_DENS_STRAT_day_mean_1992-01-02_ECCO_V4r4_latlon_0p50deg {
dimensions:
	time = 1 ;
	Z = 50 ;
	latitude = 360 ;
	longitude = 720 ;
	nv = 2 ;
variables:
	int time(time) ;
		time:axis = "T" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "center time of averaging period or time of snapshot" ;
		time:standard_name = "time" ;
		time:units = "days since 1992-01-02 12:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float Z(Z) ;
		Z:axis = "Z" ;
		Z:bounds = "Z_bnds" ;
		Z:comment = "depth at center of model grid cell.  non-uniform vertical spacing" ;
		Z:coverage_content_type = "coordinate" ;
		Z:long_name = "depth" ;
		Z:standard_name = "depth" ;
		Z:units = "m" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:comment = "uniform grid spacing from -89.75 to 89.75 by 0.5" ;
		latitude:coverage_content_type = "coordinate" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:comment = "uniform grid spacing from -179.75 to 179.75 by 0.5" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	int time_step(time) ;
		time_step:coverage_content_type = "coordinate" ;
		time_step:long_name = "model time step [hours since 1992-01-01T12:00:00" ;
		time_step:units = "hours" ;
	float RHOAnoma(time, Z, latitude, longitude) ;
		RHOAnoma:_FillValue = 9.96921e+36f ;
		RHOAnoma:comment = "In-situ seawater density anomaly relative to the reference density, rhoConst, of 1029 kg m-3.. " ;
		RHOAnoma:coverage_content_type = "modelResult" ;
		RHOAnoma:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SALINITY/DENSITY" ;
		RHOAnoma:internal\ note = "INCLUDE HFACC FOR VOLUME MEAN CALCULATIONS" ;
		RHOAnoma:long_name = "In-situ seawater density anomaly" ;
		RHOAnoma:units = "kg m-3" ;
		RHOAnoma:coordinates = "time Z latitude longitude time_step" ;
	float latitude_bnds(latitude, nv) ;
		latitude_bnds:coverage_content_type = "coordinate" ;
		latitude_bnds:long_name = "latitude bounds of lat-lon grid cells" ;
	float longitude_bnds(longitude, nv) ;
		longitude_bnds:coverage_content_type = "coordinate" ;
		longitude_bnds:long_name = "longitude bounds of lat-lon grid cells" ;
	float Z_bnds(Z, nv) ;
		Z_bnds:comment = "identical to model grid depth bounds" ;
		Z_bnds:coverage_content_type = "coordinate" ;
		Z_bnds:long_name = "depth bounds of grid cells" ;
	int time_bnds(time, nv) ;
		time_bnds:coverage_content_type = "coordinate" ;
		time_bnds:long_name = "start and stop time of period or time of snapshot" ;
		time_bnds:units = "days since 1992-01-02 00:00:00" ;
		time_bnds:calendar = "proleptic_gregorian" ;
	float DRHODR(time, Z, latitude, longitude) ;
		DRHODR:_FillValue = 9.96921e+36f ;
		DRHODR:comment = "Density stratification: d(sigma) d z-1. Note: density computations are done with in-situ density.  The vertical derivatives of in-situ density and locally-referenced potential density are identical  The equation of state is a modified UNESCO formula by Jackett and McDougall (1995), which uses the model variable potential temperature as input assuming a horizontally and temporally constant pressure of $p_0=-g \rho_{0} z$." ;
		DRHODR:coverage_content_type = "modelResult" ;
		DRHODR:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SALINITY/DENSITY" ;
		DRHODR:internal\ note = "is stratification calculated on z* or z coordinates?" ;
		DRHODR:long_name = "Density stratification" ;
		DRHODR:units = "kg m-3 m-1" ;
		DRHODR:coordinates = "time Z latitude longitude time_step" ;
	float PHIHYD(time, Z, latitude, longitude) ;
		PHIHYD:_FillValue = 9.96921e+36f ;
		PHIHYD:comment = "Anomaly of hydrostatic ocean pressure normalized by a reference density (rhoConst) with respect to gz*(k,t), where g is acceleration due to gravity, 9.81 m s-2,  z*(k,t) is model depth at level k and time t, and rhoConst is 1029 kg m-3.. Note: also referred to in some contexts as hydrostatic pressure potential anomaly.  PHIHYD is calculated with respect to the model\'s time-varying grid cell thicknesses allowed by z* coordinate system. See PHIHYDcR for hydrostatic pressure potential anomaly calculated using time-invariant grid cell thicknesses. PHIHYD is NOT corrected for spurious mass fluxes incurred by density changes in the Boussinesq volume-conserving model (Greatbatch correction) (see sterGloH). " ;
		PHIHYD:coverage_content_type = "modelResult" ;
		PHIHYD:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; OCEAN PRESSURE; WATER PRESSURE" ;
		PHIHYD:long_name = "Ocean hydrostatic pressure anomaly" ;
		PHIHYD:units = "m2 s-2" ;
		PHIHYD:coordinates = "time Z latitude longitude time_step" ;

// global attributes:
		:acknowledgement = "This research was carried out by the Jet Propulsion Laboratory, managed by the California Institute of Technology under a contract with the National Aeronautics and Space Administration." ;
		:author = "Ian Fenty and Ou Wang" ;
		:cdm_data_type = "Grid" ;
		:comment = "These fields are provided on a regular lat-lon grid. They have been mapped to the regular lat-lon grid from the original ECCO lat-lon-cap 90 (llc90) native model grid." ;
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:coordinates = "time Z latitude longitude time_step latitude_bnds longitude_bnds Z_bnds time_bnds" ;
		:creator_email = "ecco-group@mit.edu" ;
		:creator_institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:creator_name = "ECCO Consortium" ;
		:creator_type = "group" ;
		:creator_url = "https://ecco.jpl.nasa.gov" ;
		:date_created = "TBD_DATASET" ;
		:date_issued = "2020-09-02T15:32:14.761407" ;
		:date_metadata_modified = "2020-09-02T15:32:14.761405" ;
		:date_modified = "2020-09-02T15:32:14.761387" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 90. ;
		:geospatial_lat_min = -90. ;
		:geospatial_lat_resolution = 0.5 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 180. ;
		:geospatial_lon_min = -180. ;
		:geospatial_lon_resolution = 0.5 ;
		:geospatial_lon_units = "degrees_east" ;
		:grid_mapping_name = "latitude_longitude" ;
		:history = "Inaugural release of an ECCO \"Central Estimate\" solution to PO.DAAC" ;
		:id = "TBD_DOI" ;
		:institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:keywords = "ECCO, State Estimate, Estimating the Circulation and Climate of the Ocean" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "Public Domain" ;
		:naming_authority = "gov.nasa.jpl" ;
		:nx = 720 ;
		:ny = 360 ;
		:platform = "ERS-1/2, TOPEX/Poseidon, GFO, ENVISAT, Jason-1, Jason-2, CryoSat-2, SARAL/AltiKa, Jason-3, AVHRR, Aquarius, SSM/I, SSMIS, GRACE, DTU17MDT, Argo, WOCE, GO-SHIP, MEOP, ITP" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:processing_level = "L4" ;
		:product_name = "TBD_FILENAME" ;
		:product_time_coverage_end = "2017-12-31T12:00:00" ;
		:product_time_coverage_start = "1992-01-01T12:00:00" ;
		:product_version = "Version 4, Release 4" ;
		:program = "NASA Physical Oceanography, Cryosphere, Modeling, Analysis, and Prediction (MAP)" ;
		:project = "Estimating the Circulation and Climate of the Ocean (ECCO)" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_institution = "PO.DAAC" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center (PO.DAAC)" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:references = "ECCO Consortium, Fukumori, I., Wang, O., Fenty, I., Forget, G., Heimbach, P., & Ponte, R. M. 2020. Synopsis of the ECCO Central Production Global Ocean and Sea-Ice State Estimate (Version 4 Release 4).doi:10.5281/zenodo.3765929" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:summary = "ocean density, stratification, and hydrostatic pressure" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_end = "1992-01-03T00:00:00.000000000" ;
		:time_coverage_resolution = "P1D" ;
		:time_coverage_start = "1992-01-02T00:00:00.000000000" ;
		:title = "ocean density, stratification, and hydrostatic pressure" ;
		:uuid = "TBD_DATASET" ;
}
