netcdf SURFACE_HEAT_FLUXES_day_mean_1992-01-01_ECCO_V4r4_latlon_0p50deg {
dimensions:
	time = 1 ;
	latitude = 360 ;
	longitude = 720 ;
	nv = 2 ;
variables:
	int time(time) ;
		time:axis = "T" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "center time of averaging period or time of snapshot" ;
		time:standard_name = "time" ;
		time:units = "days since 1992-01-01 12:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:comment = "uniform grid spacing from -89.75 to 89.75 by 0.5" ;
		latitude:coverage_content_type = "coordinate" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:comment = "uniform grid spacing from -179.75 to 179.75 by 0.5" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	int time_step(time) ;
		time_step:coverage_content_type = "coordinate" ;
		time_step:long_name = "model time step [hours since 1992-01-01T12:00:00" ;
		time_step:units = "hours" ;
	float EXFhl(time, latitude, longitude) ;
		EXFhl:_FillValue = 9.96921e+36f ;
		EXFhl:comment = "Open ocean latent heat flux. Note: calculated from the bulk formula following Large and Yeager, 2004, NCAR/TN-460+STR." ;
		EXFhl:coverage_content_type = "modelResult" ;
		EXFhl:direction = ">0 increases potential temperature (THETA)" ;
		EXFhl:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE; OCEAN HEAT BUDGET; HEAT FLUX" ;
		EXFhl:long_name = "Air-sea latent heat flux" ;
		EXFhl:standard_name = "surface_downward_latent_heat_flux" ;
		EXFhl:units = "W m-2" ;
		EXFhl:coordinates = "time latitude longitude time_step" ;
	float latitude_bnds(latitude, nv) ;
		latitude_bnds:coverage_content_type = "coordinate" ;
		latitude_bnds:long_name = "latitude bounds of lat-lon grid cells" ;
	float longitude_bnds(longitude, nv) ;
		longitude_bnds:coverage_content_type = "coordinate" ;
		longitude_bnds:long_name = "longitude bounds of lat-lon grid cells" ;
	int time_bnds(time, nv) ;
		time_bnds:coverage_content_type = "coordinate" ;
		time_bnds:long_name = "start and stop time of period or time of snapshot" ;
		time_bnds:units = "days since 1992-01-01 00:00:00" ;
		time_bnds:calendar = "proleptic_gregorian" ;
	float EXFhs(time, latitude, longitude) ;
		EXFhs:_FillValue = 9.96921e+36f ;
		EXFhs:comment = "Open ocean sensible heat flux. Note: calculated from the bulk formula following Large and Yeager, 2004, NCAR/TN-460+STR." ;
		EXFhs:coverage_content_type = "modelResult" ;
		EXFhs:direction = ">0 increases potential temperature (THETA)" ;
		EXFhs:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE; OCEAN HEAT BUDGET; HEAT FLUX" ;
		EXFhs:long_name = "Air-sea sensible heat flux" ;
		EXFhs:standard_name = "surface_downward_sensible_heat_flux" ;
		EXFhs:units = "W m-2" ;
		EXFhs:coordinates = "time latitude longitude time_step" ;
	float EXFlwdn(time, latitude, longitude) ;
		EXFlwdn:_FillValue = 9.96921e+36f ;
		EXFlwdn:comment = "Downward longwave radiative flux. Note: sum of ERA-Interim downward longwave radiation and the control adjustment." ;
		EXFlwdn:coverage_content_type = "modelResult" ;
		EXFlwdn:direction = ">0 increases potential temperature (THETA)" ;
		EXFlwdn:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE;ATMOSPHERIC RADIATION; HEAT FLUX; LONGWAVE RADIATION; RADIATIVE FORCING; RADIATIVE FLUX" ;
		EXFlwdn:long_name = "Downward longwave radiative flux" ;
		EXFlwdn:standard_name = "surface_downwelling_longwave_flux_in_air" ;
		EXFlwdn:units = "W m-2" ;
		EXFlwdn:coordinates = "time latitude longitude time_step" ;
	float EXFswdn(time, latitude, longitude) ;
		EXFswdn:_FillValue = 9.96921e+36f ;
		EXFswdn:comment = "Downward shortwave radiative flux. Note: sum of ERA-Interim downward shortwave radiation and the control adjustment." ;
		EXFswdn:coverage_content_type = "modelResult" ;
		EXFswdn:direction = ">0 increases potential temperature (THETA)" ;
		EXFswdn:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE;ATMOSPHERIC RADIATION; OCEAN HEAT BUDGET; HEAT FLUX; INCOMING SOLAR RADIATION; SHORTWAVE RADIATION; RADIATIVE FORCING; RADIATIVE FLUX" ;
		EXFswdn:long_name = "Downwelling shortwave radiative flux" ;
		EXFswdn:standard_name = "surface_downwelling_shortwave_flux_in_air" ;
		EXFswdn:units = "W m-2" ;
		EXFswdn:coordinates = "time latitude longitude time_step" ;
	float EXFqnet(time, latitude, longitude) ;
		EXFqnet:_FillValue = 9.96921e+36f ;
		EXFqnet:comment = "Open ocean net heat flux (turbulent and radiative). Note: net upward heat flux over open water, calculated as EXFlwnet+EXFswnet-EXFlh-EXFhs." ;
		EXFqnet:coverage_content_type = "modelResult" ;
		EXFqnet:direction = ">0 increases potential temperature (THETA)" ;
		EXFqnet:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE; OCEAN HEAT BUDGET; HEAT FLUX" ;
		EXFqnet:long_name = "Net air-sea heat flux" ;
		EXFqnet:units = "W m-2" ;
		EXFqnet:coordinates = "time latitude longitude time_step" ;
	float oceQnet(time, latitude, longitude) ;
		oceQnet:_FillValue = 9.96921e+36f ;
		oceQnet:comment = "Net heat flux across the ocean surface from all processes: air-sea turbulent and radiative fluxes and turbulent and conductive fluxes between the ocean and sea-ice and snow.. Note: \'oceQnet\' does not include the change in ocean heat content due to changing ocean ocean mass (\'oceFWflx\'). Mass fluxes from evaporation, precipitation, and runoff (\'EXFempmr\') happen at the same temperature as the ocean surface temperature. Consequently, EmPmR does not change ocean surface temperature. Conversely, mass fluxes due to sea-ice thickening/thinning and snow melt in the model are assumed to happen at a fixed 0C. Consequently, mass fluxes due to phase changes between seawater and sea-ice and snow induce a heat flux when the ocean surface temperaure is not 0C. The variable \'TFLUX\' does include the change in ocean heat content due to changing ocean mass." ;
		oceQnet:coverage_content_type = "modelResult" ;
		oceQnet:direction = ">0 increases potential temperature (THETA)" ;
		oceQnet:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; ATMOSPHERE; OCEAN HEAT BUDGET; HEAT FLUX" ;
		oceQnet:long_name = "Net heat flux across the ocean surface" ;
		oceQnet:units = "W m-2" ;
		oceQnet:coordinates = "time latitude longitude time_step" ;
	float SIatmQnt(time, latitude, longitude) ;
		SIatmQnt:_FillValue = 9.96921e+36f ;
		SIatmQnt:comment = "Net heat flux to the atmosphere across open water and sea-ice or snow surfaces.. Note: for sea-ice covered regions, positive \'SIatmQnt\' may have no effect on ocean potential temperature. Does NOT include the contribution to the ocean heat content from changing mass (e.g. from \'oceFWflx\'). \'TFLUX\' includes the contribution to the ocean heat content from changing mass." ;
		SIatmQnt:coverage_content_type = "modelResult" ;
		SIatmQnt:direction = ">0 upward" ;
		SIatmQnt:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SEA ICE; SNOW/ICE; HEAT FLUX" ;
		SIatmQnt:long_name = "Upward heat flux across the lower boundary of atmosphere" ;
		SIatmQnt:standard_name = "downward_heat_flux_in_air" ;
		SIatmQnt:units = "W m-2" ;
		SIatmQnt:coordinates = "time latitude longitude time_step" ;
	float TFLUX(time, latitude, longitude) ;
		TFLUX:_FillValue = 9.96921e+36f ;
		TFLUX:comment = "The rate of change of ocean heat content due to heat fluxes across the liquid surface and the addition or removal of mass. . Note: the global area integral of \'TFLUX\' and geothermal flux (geothermalFlux.bin) matches the time-derivative of ocean heat content (J/s). Unlike oceQnet, TFLUX includes the contribution to the ocean heat content from changing ocean mass (e.g. from oceFWflx)." ;
		TFLUX:coverage_content_type = "modelResult" ;
		TFLUX:direction = ">0 increases potential temperature (THETA)" ;
		TFLUX:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; OCEAN HEAT BUDGET; HEAT FLUX" ;
		TFLUX:long_name = "Rate of change of ocean heat content per m2 accounting for mass fluxes." ;
		TFLUX:units = "W m-2" ;
		TFLUX:coordinates = "time latitude longitude time_step" ;
	float EXFswnet(time, latitude, longitude) ;
		EXFswnet:_FillValue = 9.96921e+36f ;
		EXFswnet:comment = "Open ocean net shortwave radiative flux. Note: net shortwave flux net shortwave radiation over open water calculated from downward longave shortwave over open water (EXFlwdn) and ocean surface albdeo." ;
		EXFswnet:coverage_content_type = "modelResult" ;
		EXFswnet:direction = ">0 increases potential temperature (THETA)" ;
		EXFswnet:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE;ATMOSPHERIC RADIATION; OCEAN HEAT BUDGET; HEAT FLUX; INCOMING SOLAR RADIATION; NET RADIATION; SHORTWAVE RADIATION; RADIATIVE FORCING; RADIATIVE FLUX" ;
		EXFswnet:long_name = "Net open ocean shortwave radiative flux" ;
		EXFswnet:standard_name = "surface_net_downward_shortwave_flux" ;
		EXFswnet:units = "W m-2" ;
		EXFswnet:coordinates = "time latitude longitude time_step" ;
	float EXFlwnet(time, latitude, longitude) ;
		EXFlwnet:_FillValue = 9.96921e+36f ;
		EXFlwnet:comment = "Open ocean net upward longwave radiative flux. Note: net longwave radiation over open water calculated from downward longave radiation over open water (EXFlwdn) and Stefan-Boltzman." ;
		EXFlwnet:coverage_content_type = "modelResult" ;
		EXFlwnet:direction = ">0 increases potential temperature (THETA)" ;
		EXFlwnet:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; ATMOSPHERE;ATMOSPHERIC RADIATION; OCEAN HEAT BUDGET; HEAT FLUX; LONGWAVE RADIATION; OUTGOING LONGWAVE RADIATION; NET RADIATION; RADIATIVE FORCING; RADIATIVE FLUX" ;
		EXFlwnet:long_name = "Net longwave radiative flux" ;
		EXFlwnet:standard_name = "surface_net_downward_longwave_flux" ;
		EXFlwnet:units = "W m-2" ;
		EXFlwnet:coordinates = "time latitude longitude time_step" ;
	float oceQsw(time, latitude, longitude) ;
		oceQsw:_FillValue = 9.96921e+36f ;
		oceQsw:comment = "Net shortwave radiative flux across the ocean surface. Note: Shortwave radiation penetrates below the surface grid cell." ;
		oceQsw:coverage_content_type = "modelResult" ;
		oceQsw:direction = ">0 increases potential temperature (THETA)" ;
		oceQsw:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; ATMOSPHERE;ATMOSPHERIC RADIATION; OCEAN HEAT BUDGET; HEAT FLUX; INCOMING SOLAR RADIATION; SHORTWAVE RADIATION; RADIATIVE FORCING; RADIATIVE FLUX" ;
		oceQsw:long_name = "Net shortwave radiative flux across the ocean surface" ;
		oceQsw:units = "W m-2" ;
		oceQsw:coordinates = "time latitude longitude time_step" ;
	float SIaaflux(time, latitude, longitude) ;
		SIaaflux:_FillValue = 9.96921e+36f ;
		SIaaflux:comment = "Heat flux associated with the temperature difference between sea surface temperature and sea-ice (assume 0 degree C in the model). Note: heat flux needed to melt/freeze sea-ice at 0 degC to sea water at the ocean surface (at sea surface temperature), excluding the latent heat of fusion." ;
		SIaaflux:coverage_content_type = "modelResult" ;
		SIaaflux:direction = ">0 decrease potential temperature (THETA)" ;
		SIaaflux:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; SEA ICE; SNOW/ICE; HEAT FLUX" ;
		SIaaflux:long_name = "Conservative ocean and sea-ice advective heat flux adjustment" ;
		SIaaflux:units = "W m-2" ;
		SIaaflux:coordinates = "time latitude longitude time_step" ;

// global attributes:
		:acknowledgement = "This research was carried out by the Jet Propulsion Laboratory, managed by the California Institute of Technology under a contract with the National Aeronautics and Space Administration." ;
		:author = "Ian Fenty and Ou Wang" ;
		:cdm_data_type = "Grid" ;
		:comment = "These fields are provided on a regular lat-lon grid. They have been mapped to the regular lat-lon grid from the original ECCO lat-lon-cap 90 (llc90) native model grid." ;
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:coordinates = "time latitude longitude time_step latitude_bnds longitude_bnds time_bnds" ;
		:creator_email = "ecco-group@mit.edu" ;
		:creator_institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:creator_name = "ECCO Consortium" ;
		:creator_type = "group" ;
		:creator_url = "https://ecco.jpl.nasa.gov" ;
		:date_created = "TBD_DATASET" ;
		:date_issued = "2020-09-02T15:33:17.355935" ;
		:date_metadata_modified = "2020-09-02T15:33:17.355932" ;
		:date_modified = "2020-09-02T15:33:17.355923" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 90. ;
		:geospatial_lat_min = -90. ;
		:geospatial_lat_resolution = 0.5 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 180. ;
		:geospatial_lon_min = -180. ;
		:geospatial_lon_resolution = 0.5 ;
		:geospatial_lon_units = "degrees_east" ;
		:grid_mapping_name = "latitude_longitude" ;
		:history = "Inaugural release of an ECCO \"Central Estimate\" solution to PO.DAAC" ;
		:id = "TBD_DOI" ;
		:institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:keywords = "ECCO, State Estimate, Estimating the Circulation and Climate of the Ocean" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "Public Domain" ;
		:naming_authority = "gov.nasa.jpl" ;
		:nx = 720 ;
		:ny = 360 ;
		:platform = "ERS-1/2, TOPEX/Poseidon, GFO, ENVISAT, Jason-1, Jason-2, CryoSat-2, SARAL/AltiKa, Jason-3, AVHRR, Aquarius, SSM/I, SSMIS, GRACE, DTU17MDT, Argo, WOCE, GO-SHIP, MEOP, ITP" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:processing_level = "L4" ;
		:product_name = "TBD_FILENAME" ;
		:product_time_coverage_end = "2017-12-31T12:00:00" ;
		:product_time_coverage_start = "1992-01-01T12:00:00" ;
		:product_version = "Version 4, Release 4" ;
		:program = "NASA Physical Oceanography, Cryosphere, Modeling, Analysis, and Prediction (MAP)" ;
		:project = "Estimating the Circulation and Climate of the Ocean (ECCO)" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_institution = "PO.DAAC" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center (PO.DAAC)" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:references = "ECCO Consortium, Fukumori, I., Wang, O., Fenty, I., Forget, G., Heimbach, P., & Ponte, R. M. 2020. Synopsis of the ECCO Central Production Global Ocean and Sea-Ice State Estimate (Version 4 Release 4).doi:10.5281/zenodo.3765929" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:summary = "ocean and sea-ice surface heat fluxes" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_end = "1992-01-02T00:00:00.000000000" ;
		:time_coverage_resolution = "P1D" ;
		:time_coverage_start = "1992-01-01T00:00:00.000000000" ;
		:title = "ocean and sea-ice surface heat fluxes" ;
		:uuid = "TBD_DATASET" ;
}
