netcdf OCEAN_SURFACE_STRESS_mon_mean_1992-02_ECCO_V4r4_latlon_0p50deg {
dimensions:
	time = 1 ;
	latitude = 360 ;
	longitude = 720 ;
	nv = 2 ;
variables:
	int time(time) ;
		time:axis = "T" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "center time of averaging period or time of snapshot" ;
		time:standard_name = "time" ;
		time:units = "days since 1992-02-15 12:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:comment = "uniform grid spacing from -89.75 to 89.75 by 0.5" ;
		latitude:coverage_content_type = "coordinate" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:comment = "uniform grid spacing from -179.75 to 179.75 by 0.5" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	int time_step(time) ;
		time_step:coverage_content_type = "coordinate" ;
		time_step:long_name = "model time step [hours since 1992-01-01T12:00:00" ;
		time_step:units = "hours" ;
	float EXFtaue(time, latitude, longitude) ;
		EXFtaue:_FillValue = 9.96921e+36f ;
		EXFtaue:comment = "Zonal (east-west) component of wind stress. Note: EXFtaue is the zonal wind stress applied to the ocean and sea-ice. When sea-ice is present, the total zonal stress applied to the ocean surface is NOT EXFtaue, but a combination of the wind stress in the open water fraction (EXFtaue) and a stress from sea-ice in the ice-covered fraction (see oceTAUE). EXFtaue is calculated by interpolating the model\'s x and y components of wind stress (EXFtaux and EXFtauy) to tracer cell centers and then finding the zonal component of the interpolated vectors. It is NOT recommended to use EXFtaue and EXFtaun for momentum budget calculations because interpolating EXFtaux and EXFtauy from the model grid to the lat-lon grid introduces errors. For momentum fluxes to the ocean surface see oceTAUx and oceTAUy." ;
		EXFtaue:coverage_content_type = "modelResult" ;
		EXFtaue:direction = " >0 increases eastward velocity (EVEL)" ;
		EXFtaue:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; ATMOSPHERE; WIND STRESS" ;
		EXFtaue:long_name = "Zonal (east-west) wind stress" ;
		EXFtaue:standard_name = "surface_downward_eastward_stress" ;
		EXFtaue:units = "N m-2" ;
		EXFtaue:coordinates = "time latitude longitude time_step" ;
	float latitude_bnds(latitude, nv) ;
		latitude_bnds:coverage_content_type = "coordinate" ;
		latitude_bnds:long_name = "latitude bounds of lat-lon grid cells" ;
	float longitude_bnds(longitude, nv) ;
		longitude_bnds:coverage_content_type = "coordinate" ;
		longitude_bnds:long_name = "longitude bounds of lat-lon grid cells" ;
	int time_bnds(time, nv) ;
		time_bnds:coverage_content_type = "coordinate" ;
		time_bnds:long_name = "start and stop time of period or time of snapshot" ;
		time_bnds:units = "days since 1992-02-01 00:00:00" ;
		time_bnds:calendar = "proleptic_gregorian" ;
	float EXFtaun(time, latitude, longitude) ;
		EXFtaun:_FillValue = 9.96921e+36f ;
		EXFtaun:comment = "Meridional (north-south) component of wind stress. Note: EXFtaun is the stress applied to the ocean and sea-ice. When sea-ice is present, the total meridional stress applied to the ocean surface is NOT EXFtaun, but a combination of the wind stress in the open water fraction (EXFtaun) and a stress from sea-ice in the ice-covered fraction (see oceTAUN).  EXFtaun is calculated by interpolating the model\'s x and y components of wind stress (EXFtaux and EXFtauy) to tracer cell centers and then determining the meridional component of the interpolated vectors. It is NOT recommended to use EXFtaue and EXFtaun for momentum budget calculations because interpolating EXFtaux and EXFtauy from the model grid to the lat-lon grid introduces errors. For momentum fluxes to the ocean surface see oceTAUx and oceTAUy." ;
		EXFtaun:coverage_content_type = "modelResult" ;
		EXFtaun:direction = " >0 increases northward velocity (NVEL)" ;
		EXFtaun:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; ATMOSPHERE; WIND STRESS" ;
		EXFtaun:long_name = "Meridional (north-south) wind stress" ;
		EXFtaun:standard_name = "surface_downward_northward_stress" ;
		EXFtaun:units = "N m-2" ;
		EXFtaun:coordinates = "time latitude longitude time_step" ;
	float oceTAUE(time, latitude, longitude) ;
		oceTAUE:_FillValue = 9.96921e+36f ;
		oceTAUE:comment = "Zonal (east-west) component of ocean surface stress due to wind and sea-ice. Note: oceTAUE is calculated by interpolating the model\'s x and y components of ocean surface stress (oceTAUX and oceTAUY) to tracer cell centers and then finding the zonal component of the interpolated vectors." ;
		oceTAUE:coverage_content_type = "modelResult" ;
		oceTAUE:direction = " >0 increases eastward velocity (EVEL)" ;
		oceTAUE:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; ATMOSPHERE; WIND STRESS" ;
		oceTAUE:long_name = "Zonal (east-west) ocean surface stress" ;
		oceTAUE:standard_name = "surface_downward_eastward_stress" ;
		oceTAUE:units = "N m-2" ;
		oceTAUE:coordinates = "time latitude longitude time_step" ;
	float oceTAUN(time, latitude, longitude) ;
		oceTAUN:_FillValue = 9.96921e+36f ;
		oceTAUN:comment = "Meridional (north-south) component of ocean surface stress due to wind and sea-ice. Note: oceTAUN is calculated by interpolating the model\'s x and y components of ocean surface stress (oceTAUX and oceTAUY) to tracer cell centers and then finding the meridional component of the interpolated vectors." ;
		oceTAUN:coverage_content_type = "modelResult" ;
		oceTAUN:direction = " >0 increases northward velocity (NVEL)" ;
		oceTAUN:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; ATMOSPHERE; WIND STRESS" ;
		oceTAUN:long_name = "Meridional (north-south) ocean surface stress" ;
		oceTAUN:standard_name = "surface_downward_northward_stress" ;
		oceTAUN:units = "N m-2" ;
		oceTAUN:coordinates = "time latitude longitude time_step" ;

// global attributes:
		:acknowledgement = "This research was carried out by the Jet Propulsion Laboratory, managed by the California Institute of Technology under a contract with the National Aeronautics and Space Administration." ;
		:author = "Ian Fenty and Ou Wang" ;
		:cdm_data_type = "Grid" ;
		:comment = "These fields are provided on a regular lat-lon grid. They have been mapped to the regular lat-lon grid from the original ECCO lat-lon-cap 90 (llc90) native model grid." ;
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:coordinates = "time latitude longitude time_step latitude_bnds longitude_bnds time_bnds" ;
		:creator_email = "ecco-group@mit.edu" ;
		:creator_institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:creator_name = "ECCO Consortium" ;
		:creator_type = "group" ;
		:creator_url = "https://ecco.jpl.nasa.gov" ;
		:date_created = "TBD_DATASET" ;
		:date_issued = "2020-09-02T15:35:18.483841" ;
		:date_metadata_modified = "2020-09-02T15:35:18.483838" ;
		:date_modified = "2020-09-02T15:35:18.483827" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 90. ;
		:geospatial_lat_min = -90. ;
		:geospatial_lat_resolution = 0.5 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 180. ;
		:geospatial_lon_min = -180. ;
		:geospatial_lon_resolution = 0.5 ;
		:geospatial_lon_units = "degrees_east" ;
		:grid_mapping_name = "latitude_longitude" ;
		:history = "Inaugural release of an ECCO \"Central Estimate\" solution to PO.DAAC" ;
		:id = "TBD_DOI" ;
		:institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:keywords = "ECCO, State Estimate, Estimating the Circulation and Climate of the Ocean" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "Public Domain" ;
		:naming_authority = "gov.nasa.jpl" ;
		:nx = 720 ;
		:ny = 360 ;
		:platform = "ERS-1/2, TOPEX/Poseidon, GFO, ENVISAT, Jason-1, Jason-2, CryoSat-2, SARAL/AltiKa, Jason-3, AVHRR, Aquarius, SSM/I, SSMIS, GRACE, DTU17MDT, Argo, WOCE, GO-SHIP, MEOP, ITP" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:processing_level = "L4" ;
		:product_name = "TBD_FILENAME" ;
		:product_time_coverage_end = "2017-12-31T12:00:00" ;
		:product_time_coverage_start = "1992-01-01T12:00:00" ;
		:product_version = "Version 4, Release 4" ;
		:program = "NASA Physical Oceanography, Cryosphere, Modeling, Analysis, and Prediction (MAP)" ;
		:project = "Estimating the Circulation and Climate of the Ocean (ECCO)" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_institution = "PO.DAAC" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center (PO.DAAC)" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:references = "ECCO Consortium, Fukumori, I., Wang, O., Fenty, I., Forget, G., Heimbach, P., & Ponte, R. M. 2020. Synopsis of the ECCO Central Production Global Ocean and Sea-Ice State Estimate (Version 4 Release 4).doi:10.5281/zenodo.3765929" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:summary = "ocean surface stress over open water fraction (EXF*) and total over open water and ice-covered fractions (oceTAU*) " ;
		:time_coverage_duration = "P1M" ;
		:time_coverage_end = "1992-03-01T00:00:00.000000000" ;
		:time_coverage_resolution = "P1M" ;
		:time_coverage_start = "1992-02-01T00:00:00.000000000" ;
		:title = "ocean surface stress" ;
		:uuid = "TBD_DATASET" ;
}
