netcdf MIXED_LAYER_DEPTH_mon_mean_1992-02_ECCO_V4r4_latlon_0p50deg {
dimensions:
	time = 1 ;
	latitude = 360 ;
	longitude = 720 ;
	nv = 2 ;
variables:
	int time(time) ;
		time:axis = "T" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "center time of averaging period or time of snapshot" ;
		time:standard_name = "time" ;
		time:units = "days since 1992-02-15 12:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:comment = "uniform grid spacing from -89.75 to 89.75 by 0.5" ;
		latitude:coverage_content_type = "coordinate" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:comment = "uniform grid spacing from -179.75 to 179.75 by 0.5" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	int time_step(time) ;
		time_step:coverage_content_type = "coordinate" ;
		time_step:long_name = "model time step [hours since 1992-01-01T12:00:00" ;
		time_step:units = "hours" ;
	float MXLDEPTH(time, latitude, longitude) ;
		MXLDEPTH:_FillValue = 9.96921e+36f ;
		MXLDEPTH:comment = "Mixed-layer depth as determined by the depth where waters are first 0.8 degrees Celsius colder than the surface. See Kara et al. (JGR, 2000). . Note: the Kara et al. criterion may not be appropriate for some applications.  If needed, mixed layer depth can be calculated using different criteria. See vertical density stratification (DRHODR) and density anomaly (RHOAnoma)." ;
		MXLDEPTH:coverage_content_type = "modelResult" ;
		MXLDEPTH:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS; OCEAN MIXED LAYER" ;
		MXLDEPTH:long_name = "Mixed-layer depth diagnosed using the temperature difference criterion of Kara et al., 2000" ;
		MXLDEPTH:standard_name = "ocean_mixed_layer_thickness" ;
		MXLDEPTH:units = "m" ;
		MXLDEPTH:coordinates = "time latitude longitude time_step" ;
	float latitude_bnds(latitude, nv) ;
		latitude_bnds:coverage_content_type = "coordinate" ;
		latitude_bnds:long_name = "latitude bounds of lat-lon grid cells" ;
	float longitude_bnds(longitude, nv) ;
		longitude_bnds:coverage_content_type = "coordinate" ;
		longitude_bnds:long_name = "longitude bounds of lat-lon grid cells" ;
	int time_bnds(time, nv) ;
		time_bnds:coverage_content_type = "coordinate" ;
		time_bnds:long_name = "start and stop time of period or time of snapshot" ;
		time_bnds:units = "days since 1992-02-01 00:00:00" ;
		time_bnds:calendar = "proleptic_gregorian" ;

// global attributes:
		:acknowledgement = "This research was carried out by the Jet Propulsion Laboratory, managed by the California Institute of Technology under a contract with the National Aeronautics and Space Administration." ;
		:author = "Ian Fenty and Ou Wang" ;
		:cdm_data_type = "Grid" ;
		:comment = "These fields are provided on a regular lat-lon grid. They have been mapped to the regular lat-lon grid from the original ECCO lat-lon-cap 90 (llc90) native model grid." ;
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:coordinates = "time latitude longitude time_step latitude_bnds longitude_bnds time_bnds" ;
		:creator_email = "ecco-group@mit.edu" ;
		:creator_institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:creator_name = "ECCO Consortium" ;
		:creator_type = "group" ;
		:creator_url = "https://ecco.jpl.nasa.gov" ;
		:date_created = "TBD_DATASET" ;
		:date_issued = "2020-09-02T15:35:15.244365" ;
		:date_metadata_modified = "2020-09-02T15:35:15.244363" ;
		:date_modified = "2020-09-02T15:35:15.244354" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 90. ;
		:geospatial_lat_min = -90. ;
		:geospatial_lat_resolution = 0.5 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 180. ;
		:geospatial_lon_min = -180. ;
		:geospatial_lon_resolution = 0.5 ;
		:geospatial_lon_units = "degrees_east" ;
		:grid_mapping_name = "latitude_longitude" ;
		:history = "Inaugural release of an ECCO \"Central Estimate\" solution to PO.DAAC" ;
		:id = "TBD_DOI" ;
		:institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:keywords = "ECCO, State Estimate, Estimating the Circulation and Climate of the Ocean" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "Public Domain" ;
		:naming_authority = "gov.nasa.jpl" ;
		:nx = 720 ;
		:ny = 360 ;
		:platform = "ERS-1/2, TOPEX/Poseidon, GFO, ENVISAT, Jason-1, Jason-2, CryoSat-2, SARAL/AltiKa, Jason-3, AVHRR, Aquarius, SSM/I, SSMIS, GRACE, DTU17MDT, Argo, WOCE, GO-SHIP, MEOP, ITP" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:processing_level = "L4" ;
		:product_name = "TBD_FILENAME" ;
		:product_time_coverage_end = "2017-12-31T12:00:00" ;
		:product_time_coverage_start = "1992-01-01T12:00:00" ;
		:product_version = "Version 4, Release 4" ;
		:program = "NASA Physical Oceanography, Cryosphere, Modeling, Analysis, and Prediction (MAP)" ;
		:project = "Estimating the Circulation and Climate of the Ocean (ECCO)" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_institution = "PO.DAAC" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center (PO.DAAC)" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:references = "ECCO Consortium, Fukumori, I., Wang, O., Fenty, I., Forget, G., Heimbach, P., & Ponte, R. M. 2020. Synopsis of the ECCO Central Production Global Ocean and Sea-Ice State Estimate (Version 4 Release 4).doi:10.5281/zenodo.3765929" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:summary = "mixed layer depth" ;
		:time_coverage_duration = "P1M" ;
		:time_coverage_end = "1992-03-01T00:00:00.000000000" ;
		:time_coverage_resolution = "P1M" ;
		:time_coverage_start = "1992-02-01T00:00:00.000000000" ;
		:title = "mixed layer depth" ;
		:uuid = "TBD_DATASET" ;
}
