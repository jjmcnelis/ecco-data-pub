netcdf GM_OCEAN_BOLUS_VELOCITY_day_mean_1992-01-01_ECCO_V4r4_latlon_0p50deg {
dimensions:
	time = 1 ;
	Z = 50 ;
	latitude = 360 ;
	longitude = 720 ;
	nv = 2 ;
variables:
	int time(time) ;
		time:axis = "T" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "center time of averaging period or time of snapshot" ;
		time:standard_name = "time" ;
		time:units = "days since 1992-01-01 12:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float Z(Z) ;
		Z:axis = "Z" ;
		Z:bounds = "Z_bnds" ;
		Z:comment = "depth at center of model grid cell.  non-uniform vertical spacing" ;
		Z:coverage_content_type = "coordinate" ;
		Z:long_name = "depth" ;
		Z:standard_name = "depth" ;
		Z:units = "m" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:comment = "uniform grid spacing from -89.75 to 89.75 by 0.5" ;
		latitude:coverage_content_type = "coordinate" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:comment = "uniform grid spacing from -179.75 to 179.75 by 0.5" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	int time_step(time) ;
		time_step:coverage_content_type = "coordinate" ;
		time_step:long_name = "model time step [hours since 1992-01-01T12:00:00" ;
		time_step:units = "hours" ;
	float EVELSTAR(time, Z, latitude, longitude) ;
		EVELSTAR:_FillValue = 9.96921e+36f ;
		EVELSTAR:comment = "Zonal (east-west) component of the Gent-McWilliams bolus ocean velocity. Note: EVELSTAR is calculated by interpolating the model\'s x and y components of GM bolus ocean velocity (UVELSTAR and VVELSTAR) to tracer cell centers and then finding the zonal components of the interpolated vectors. One should take care when interpreting bolus velocities interpolated from the ECCO native model grid because interpolating from the model grid to the lat-lon grid introduces errors. Some closed buget calculations require bolus velocity terms on the native model grid." ;
		EVELSTAR:coverage_content_type = "modelResult" ;
		EVELSTAR:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS;OCEAN CURRENTS; OCEAN CIRCULATION" ;
		EVELSTAR:long_name = "Gent-McWilliams zonal (east-west) bolus velocity" ;
		EVELSTAR:standard_name = "eastward_sea_water_velocity_due_to_parameterized_mesoscale_eddies" ;
		EVELSTAR:units = "m s-1" ;
		EVELSTAR:coordinates = "time Z latitude longitude time_step" ;
	float latitude_bnds(latitude, nv) ;
		latitude_bnds:coverage_content_type = "coordinate" ;
		latitude_bnds:long_name = "latitude bounds of lat-lon grid cells" ;
	float longitude_bnds(longitude, nv) ;
		longitude_bnds:coverage_content_type = "coordinate" ;
		longitude_bnds:long_name = "longitude bounds of lat-lon grid cells" ;
	float Z_bnds(Z, nv) ;
		Z_bnds:comment = "identical to model grid depth bounds" ;
		Z_bnds:coverage_content_type = "coordinate" ;
		Z_bnds:long_name = "depth bounds of grid cells" ;
	int time_bnds(time, nv) ;
		time_bnds:coverage_content_type = "coordinate" ;
		time_bnds:long_name = "start and stop time of period or time of snapshot" ;
		time_bnds:units = "days since 1992-01-01 00:00:00" ;
		time_bnds:calendar = "proleptic_gregorian" ;
	float NVELSTAR(time, Z, latitude, longitude) ;
		NVELSTAR:_FillValue = 9.96921e+36f ;
		NVELSTAR:comment = "Meridional (north-south) component of the Gent-McWilliams bolus ocean velocity. Note: NVELSTAR is calculated by interpolating the model\'s x and y components of GM bolus ocean velocity (UVELSTAR and VVELSTAR) to tracer cell centers and then finding the meridional components of the interpolated vectors.  One should take care when interpreting bolus velocities interpolated from the ECCO native model grid because interpolating from the model grid to the lat-lon grid introduces errors. Some closed buget calculations require bolus velocity terms on the native model grid" ;
		NVELSTAR:coverage_content_type = "modelResult" ;
		NVELSTAR:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS;OCEAN CURRENTS; OCEAN CIRCULATION" ;
		NVELSTAR:long_name = "Gent-McWilliams meridional (north-south) bolus velocity" ;
		NVELSTAR:standard_name = "northward_sea_water_velocity_due_to_parameterized_mesoscale_eddies" ;
		NVELSTAR:units = "m s-1" ;
		NVELSTAR:coordinates = "time Z latitude longitude time_step" ;
	float WVELSTAR(time, Z, latitude, longitude) ;
		WVELSTAR:_FillValue = 9.96921e+36f ;
		WVELSTAR:comment = "Vertical component of the Gent-McWilliams bolus ocean velocity. Note: in the Arakawa-C grid used in ECCO, vertical velocities are staggered relative to the tracer cell centers with values at the TOP and BOTTOM faces of each grid cell." ;
		WVELSTAR:coverage_content_type = "modelResult" ;
		WVELSTAR:gmcd_keywords = "REANALYSIS MODELS; EARTH SCIENCE; GCM; OCEANS;OCEAN CURRENTS; OCEAN CIRCULATION" ;
		WVELSTAR:long_name = "Gent-McWilliams vertical bolus velocity" ;
		WVELSTAR:standard_name = "upward_sea_water_velocity_due_to_parameterized_mesoscale_eddies" ;
		WVELSTAR:units = "m s-1" ;
		WVELSTAR:coordinates = "time Z latitude longitude time_step" ;

// global attributes:
		:acknowledgement = "This research was carried out by the Jet Propulsion Laboratory, managed by the California Institute of Technology under a contract with the National Aeronautics and Space Administration." ;
		:author = "Ian Fenty and Ou Wang" ;
		:cdm_data_type = "Grid" ;
		:comment = "These fields are provided on a regular lat-lon grid. They have been mapped to the regular lat-lon grid from the original ECCO lat-lon-cap 90 (llc90) native model grid." ;
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:coordinates = "time Z latitude longitude time_step latitude_bnds longitude_bnds Z_bnds time_bnds" ;
		:creator_email = "ecco-group@mit.edu" ;
		:creator_institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:creator_name = "ECCO Consortium" ;
		:creator_type = "group" ;
		:creator_url = "https://ecco.jpl.nasa.gov" ;
		:date_created = "TBD_DATASET" ;
		:date_issued = "2020-09-02T15:32:55.330470" ;
		:date_metadata_modified = "2020-09-02T15:32:55.330468" ;
		:date_modified = "2020-09-02T15:32:55.330457" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 90. ;
		:geospatial_lat_min = -90. ;
		:geospatial_lat_resolution = 0.5 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 180. ;
		:geospatial_lon_min = -180. ;
		:geospatial_lon_resolution = 0.5 ;
		:geospatial_lon_units = "degrees_east" ;
		:grid_mapping_name = "latitude_longitude" ;
		:history = "Inaugural release of an ECCO \"Central Estimate\" solution to PO.DAAC" ;
		:id = "TBD_DOI" ;
		:institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:keywords = "ECCO, State Estimate, Estimating the Circulation and Climate of the Ocean" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "Public Domain" ;
		:naming_authority = "gov.nasa.jpl" ;
		:nx = 720 ;
		:ny = 360 ;
		:platform = "ERS-1/2, TOPEX/Poseidon, GFO, ENVISAT, Jason-1, Jason-2, CryoSat-2, SARAL/AltiKa, Jason-3, AVHRR, Aquarius, SSM/I, SSMIS, GRACE, DTU17MDT, Argo, WOCE, GO-SHIP, MEOP, ITP" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:processing_level = "L4" ;
		:product_name = "TBD_FILENAME" ;
		:product_time_coverage_end = "2017-12-31T12:00:00" ;
		:product_time_coverage_start = "1992-01-01T12:00:00" ;
		:product_version = "Version 4, Release 4" ;
		:program = "NASA Physical Oceanography, Cryosphere, Modeling, Analysis, and Prediction (MAP)" ;
		:project = "Estimating the Circulation and Climate of the Ocean (ECCO)" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_institution = "PO.DAAC" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center (PO.DAAC)" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:references = "ECCO Consortium, Fukumori, I., Wang, O., Fenty, I., Forget, G., Heimbach, P., & Ponte, R. M. 2020. Synopsis of the ECCO Central Production Global Ocean and Sea-Ice State Estimate (Version 4 Release 4).doi:10.5281/zenodo.3765929" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:summary = "Gent-McWilliams ocean bolus velocity" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_end = "1992-01-02T00:00:00.000000000" ;
		:time_coverage_resolution = "P1D" ;
		:time_coverage_start = "1992-01-01T00:00:00.000000000" ;
		:title = "Gent-McWilliams ocean bolus velocity" ;
		:uuid = "TBD_DATASET" ;
}
