netcdf MIXED_LAYER_DEPTH_day_mean_1992-01-02_ECCO_V4r4_latlon_0p50deg {
dimensions:
	time = 1 ;
	latitude = 360 ;
	longitude = 720 ;
	nv = 2 ;
variables:
	int time(time) ;
		time:axis = "T" ;
		time:coverage_content_type = "coordinate" ;
		time:long_name = "center time of averaging period or time of snapshot" ;
		time:standard_name = "time" ;
		time:units = "days since 1992-01-02 12:00:00" ;
		time:calendar = "proleptic_gregorian" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:comment = "uniform grid spacing from -89.75 to 89.75 by 0.5" ;
		latitude:coverage_content_type = "coordinate" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:comment = "uniform grid spacing from -179.75 to 179.75 by 0.5" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	int time_step(time) ;
		time_step:coverage_content_type = "coordinate" ;
		time_step:long_name = "model time step [hours since 1992-01-01T12:00:00]" ;
		time_step:units = "hours" ;
	float MXLDEPTH(time, latitude, longitude) ;
		MXLDEPTH:_FillValue = 9.96921e+36f ;
		MXLDEPTH:comment = "Mixed-layer depth as determined by the depth where waters are first 0.8 degrees Celsius colder than the surface. See Kara et al. (JGR, 2000). . Note: the Kara et al. criterion may not be appropriate for some applications.  If needed, mixed layer depth can be calculated using different criteria. See vertical density stratification (DRHODR) and density anomaly (RHOAnoma)." ;
		MXLDEPTH:coverage_content_type = "modelResult" ;
		MXLDEPTH:long_name = "Mixed-layer depth diagnosed using the temperature difference criterion of Kara et al., 2000" ;
		MXLDEPTH:standard_name = "ocean_mixed_layer_thickness" ;
		MXLDEPTH:units = "m" ;
		MXLDEPTH:coordinates = "time latitude longitude" ;
	float latitude_bnds(latitude, nv) ;
		latitude_bnds:coverage_content_type = "coordinate" ;
		latitude_bnds:long_name = "latitude bounds of lat-lon grid cells" ;
	float longitude_bnds(longitude, nv) ;
		longitude_bnds:coverage_content_type = "coordinate" ;
		longitude_bnds:long_name = "longitude bounds of lat-lon grid cells" ;
	int time_bnds(time, nv) ;
		time_bnds:coverage_content_type = "coordinate" ;
		time_bnds:long_name = "start and stop time of period or time of snapshot" ;
		time_bnds:units = "days since 1992-01-02 00:00:00" ;
		time_bnds:calendar = "proleptic_gregorian" ;

// global attributes:
		:acknowledgement = "This research was carried out by the Jet Propulsion Laboratory, managed by the California Institute of Technology under a contract with the National Aeronautics and Space Administration." ;
		:author = "Ian Fenty and Ou Wang" ;
		:cdm_data_type = "Grid" ;
		:comment = "These fields are provided on a regular lat-lon grid. They have been mapped to the regular lat-lon grid from the original ECCO lat-lon-cap 90 (llc90) native model grid." ;
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:creator_email = "ecco-group@mit.edu" ;
		:creator_institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:creator_name = "ECCO Consortium" ;
		:creator_type = "group" ;
		:creator_url = "https://ecco.jpl.nasa.gov" ;
		:date_created = "2020-09-03T04:19:21" ;
		:date_issued = "2020-09-03T04:19:21" ;
		:date_metadata_modified = "2020-09-03T04:19:21" ;
		:date_modified = "2020-09-03T04:19:21" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_max = 90. ;
		:geospatial_lat_min = -90. ;
		:geospatial_lat_resolution = 0.5 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 180. ;
		:geospatial_lon_min = -180. ;
		:geospatial_lon_resolution = 0.5 ;
		:geospatial_lon_units = "degrees_east" ;
		:history = "Inaugural release of an ECCO \"Central Estimate\" solution to PO.DAAC" ;
		:id = "10.5067/ECG5D-OML44" ;
		:institution = "NASA Jet Propulsion Laboratory (JPL)" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:keywords = "EARTH SCIENCE > OCEANS > OCEAN CIRCULATION > OCEAN MIXED LAYER, ECCO, State Estimate, Estimating the Circulation and Climate of the Ocean" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "Public Domain" ;
		:metadata_link = "https://cmr.earthdata.nasa.gov/search/collections.umm_json?ShortName=ECCO_L4_MIXED_LAYER_DEPTH_05DEG_DAILY_V4R4" ;
		:naming_authority = "gov.nasa.jpl" ;
		:platform = "ERS-1/2, TOPEX/Poseidon, GFO, ENVISAT, Jason-1, Jason-2, CryoSat-2, SARAL/AltiKa, Jason-3, AVHRR, Aquarius, SSM/I, SSMIS, GRACE, DTU17MDT, Argo, WOCE, GO-SHIP, MEOP, ITP" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:processing_level = "L4" ;
		:product_name = "MIXED_LAYER_DEPTH_day_mean_1992-01-02_ECCO_V4r4_latlon_0p50deg.nc" ;
		:product_time_coverage_end = "2017-12-31T12:00:00" ;
		:product_time_coverage_start = "1992-01-01T12:00:00" ;
		:product_version = "Version 4, Release 4" ;
		:program = "NASA Physical Oceanography, Cryosphere, Modeling, Analysis, and Prediction (MAP)" ;
		:project = "Estimating the Circulation and Climate of the Ocean (ECCO)" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_institution = "PO.DAAC" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center (PO.DAAC)" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:references = "ECCO Consortium, Fukumori, I., Wang, O., Fenty, I., Forget, G., Heimbach, P., & Ponte, R. M. 2020. Synopsis of the ECCO Central Production Global Ocean and Sea-Ice State Estimate (Version 4 Release 4).doi:10.5281/zenodo.3765929" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		string :summary = "This dataset provides daily average ocean mixed layer depth interpolated to a regular 0.5-degree grid as one component of a suite of ocean state estimates computed in ECCO Version 4 revision 4. \"Estimating the Circulation and Climate of the Ocean\" (ECCO) is a data assimilating model that produces optimized estimates of ocean state and flux. ECCO Version 4 release 4 (V4r4) constrains a global circulation model (MITgcm^) with diverse datasets that include satellite altimetry products like sea surface height (SSH); data derived from observations of earth’s gravity field like ocean bottom pressure (OBP); observations from diverse in situ sources like Argo, CTD, XBT, ITP, APB, Glider, and TAO mooring temperature and salinity; and numerous other datasets. ECCO V4r4 is the first of the model’s multi-decadal ocean state estimates to cover the Arctic Ocean and provide truly global coverage. It’s also the first to assimilate observations from GRACE (ocean bottom pressure) and Aquarius (sea surface salinity), and the first covering 2016 and 2017. This release represents the 25 year period from 1992 to 2017." ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_end = "1992-01-03T00:00:00" ;
		:time_coverage_resolution = "P1D" ;
		:time_coverage_start = "1992-01-02T00:00:00" ;
		:title = "ECCO Ocean Mixed Layer Depth - Daily Mean 0.5 Degree (Version 4 release 4)" ;
		:coordinates = "longitude_bnds time_step latitude_bnds time_bnds" ;
}
